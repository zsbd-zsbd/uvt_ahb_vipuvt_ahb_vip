uvt_ahb_trans.sv
